`include "ref.svh"
module imem (
    input logic [7:0] id,
    output instruction_t instr
);
    
    logic [0:255][31:0]imem;
    always_comb begin
        instr = '0;
        for (int i = 0; i < 256; i++) begin
            if (id == i) begin
                instr = imem[i];
            end            
        end
    end
    
    
    assign imem = {
        32'h00a24183,
        32'h00be0503,
        32'h017aa4aa,
        32'h00222a20,
        32'h03c5d526,
        32'h0208c100,
        32'h017f6280,
        32'h006bb582,
        32'h00e43ea4,
        32'h025b7d25,
        32'h00ebcaa2,
        32'h11cca500,
        32'h0172bea2,
        32'h03b88783,
        32'h032d2127,
        32'h0376e003,
        32'h02d45427,
        32'h038d69a0,
        32'h0192dba2,
        32'h03aaa4a2,
        32'h14b4de00,
        32'h031a9da5,
        32'h02703e22,
        32'h01864e20,
        32'h01e30083,
        32'h8f3ef280,
        32'h14fb9780,
        32'h138e6e80,
        32'h0380252f,
        32'h03a98282,
        32'h0379f3a0,
        32'h009764aa,
        32'h0001e883,
        32'h02b8542a,
        32'h0019cfa6,
        32'h01467100,
        32'h014425aa,
        32'h01a8a825,
        32'h162b2280,
        32'h033f7ea4,
        32'h02a66783,
        32'h11819400,
        32'h01787ea4,
        32'h00842827,
        32'h01c08c27,
        32'h03173226,
        32'h025daba6,
        32'h01fd3680,
        32'h00289b03,
        32'h03d70a2f,
        32'h02ada8aa,
        32'h007d2ca6,
        32'h0099f3a7,
        32'had5b9b00,
        32'h02a2a383,
        32'h017bfb00,
        32'h0102bb24,
        32'h00efc7a4,
        32'h142d4500,
        32'h009f7702,
        32'h01c6f7a0,
        32'h00212fa7,
        32'h104ed100,
        32'h01d3c7a7,
        32'h09558400,
        32'h01ef5582,
        32'h017f0127,
        32'h024b1627,
        32'h032608a4,
        32'h00c3b2a6,
        32'h0378bb83,
        32'h169b5180,
        32'h02b6d2a5,
        32'h005d2683,
        32'h14d62480,
        32'h0360a02f,
        32'h02150020,
        32'h084c3300,
        32'h03db0327,
        32'h02b439af,
        32'h02a98d24,
        32'h00c03082,
        32'h01d148a7,
        32'h02db6da5,
        32'h0807b680,
        32'h0170a402,
        32'h010f6aa7,
        32'h01194220,
        32'h01f8b322,
        32'h012ce326,
        32'h0384aa26,
        32'h00856b2a,
        32'h168fad80,
        32'h11095900,
        32'h01f72e83,
        32'h01ea33a0,
        32'h03640e2a,
        32'h0143a327,
        32'h01ab57a0,
        32'h030f7100,
        32'h0067eaaf,
        32'h03ebc6a5,
        32'h0314fba0,
        32'h02884424,
        32'h0b280480,
        32'h0046c525,
        32'h013c532f,
        32'h00c90722,
        32'h01a6c683,
        32'h03759a00,
        32'h01252c20,
        32'h02cd7caf,
        32'h03504820,
        32'h01b5ec24,
        32'h03457eaa,
        32'h035f2026,
        32'h00427780,
        32'h03feed25,
        32'h037e1825,
        32'h02c59100,
        32'h00e2bb83,
        32'h09453600,
        32'h00c3d683,
        32'h01dfa826,
        32'h0046f980,
        32'h01384ca2,
        32'h8c161500,
        32'h0088ae27,
        32'h00c374a7,
        32'h03b781af,
        32'h03ef9025,
        32'h03335203,
        32'h0229b582,
        32'h00968aa0,
        32'h02937302,
        32'h01a8172a,
        32'h12226d80,
        32'h03beae22,
        32'h005713a0,
        32'h00da9826,
        32'h02912aa2,
        32'h038efd22,
        32'h021d2326,
        32'h037405a7,
        32'h02f6d5a5,
        32'h00c87925,
        32'h03befba0,
        32'h028f84aa,
        32'h0362f4a6,
        32'h00b3e602,
        32'h013f75a7,
        32'h0028bc03,
        32'h0236a6a4,
        32'h014feea7,
        32'h0328b12a,
        32'h00106200,
        32'h03e83fa0,
        32'h02494922,
        32'h03450b03,
        32'h0065c32f,
        32'h0061c3a4,
        32'h0bfa9500,
        32'h0031f3af,
        32'h019024a5,
        32'had299c80,
        32'h01564126,
        32'h03e0ce03,
        32'h02f98802,
        32'h005c2b24,
        32'h02d300a5,
        32'h01b48a03,
        32'h013929af,
        32'h03e9d883,
        32'h8cd4d200,
        32'h01c704a4,
        32'h02196ea5,
        32'h033632a5,
        32'h02745c22,
        32'h00dcb622,
        32'h10925680,
        32'h01cc71af,
        32'h01ff9a22,
        32'h01e4e2aa,
        32'h00ced7a4,
        32'h8e200e80,
        32'h02317aa5,
        32'h03c57e20,
        32'h02338580,
        32'h00d696a5,
        32'h01714726,
        32'h00d0f5a4,
        32'h03cbf325,
        32'h011f1c83,
        32'h8ef6c180,
        32'h004f6a25,
        32'h02936824,
        32'h03ecb5a7,
        32'h038bc920,
        32'h03d831a0,
        32'h000ef6a5,
        32'h03c5ef25,
        32'h002a9da7,
        32'h038b44af,
        32'h021b5fa5,
        32'h03b45aa4,
        32'h0155eaa6,
        32'h0199bf2a,
        32'h08e69b80,
        32'h026627a5,
        32'h01bac903,
        32'h013f5682,
        32'h019da802,
        32'h028f882a,
        32'h01c93a26,
        32'h001401af,
        32'h02f19e2f,
        32'h018f38a5,
        32'h007b55a5,
        32'h0048f3af,
        32'h01258b00,
        32'h02681ea5,
        32'h022f1aa0,
        32'h13cd4480,
        32'h035d9e2f,
        32'h031bd6af,
        32'h01acaa83,
        32'h00b5cea7,
        32'h036ab4af,
        32'h037efaa6,
        32'h001bf6a5,
        32'h035c4103,
        32'h034e0020,
        32'h01559b83,
        32'h000440a2,
        32'h0a6e5b00,
        32'h08a0c000,
        32'h8f43fc00,
        32'h019f88a7,
        32'h039cea26,
        32'h00b196a5,
        32'h018a6903,
        32'h018c4300,
        32'h02ee0226,
        32'h00843a00,
        32'h02be68a0,
        32'h024849a0,
        32'h0127cd24,
        32'h03b98702,
        32'h001fcaa2,
        32'h008bca24,
        32'h00664022,
        32'h0170462f,
        32'h02d93ca2,
        32'h0316f880,
        32'h00e1bf22,
        32'h03132f00
    };
endmodule